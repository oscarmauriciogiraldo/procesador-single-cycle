module Sum1(
    input [63:0] PC,
    output [63:0] out_Sum1
    );

 assign out_Sum1 = PC + 4;


endmodule